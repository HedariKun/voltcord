module voltcord

struct Message {
pub:
	id string
	channel_id string
	guild_id string
	//author
	content string
}
